module vRAM(input 




);


logic [3:0][7:0] regs[601];




endmodule 